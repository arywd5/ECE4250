library IEEE;
use std_logic_1164.all;

entity xorGate is 
	port( x, y: in bit;
			z: out bit);
 end xorGate;	
